module contador ( 
	clk,
	clr,
	lb,
	eb,
	ec,
	display
	) ;

input  clk;
input  clr;
input  lb;
input  eb;
input  ec;
inout [6:0] display;
