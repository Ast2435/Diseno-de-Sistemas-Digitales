module registro ( 
	dato,
	clk,
	clr,
	ini,
	a0,
	lb,
	eb,
	ec
	) ;

input [5:0] dato;
input  clk;
input  clr;
input  ini;
inout [5:0] a0;
inout  lb;
inout  eb;
inout  ec;
